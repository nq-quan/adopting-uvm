//-*-
 verilog-indent-level: 3; indent-tabs-mode: nil; tab-width: 1 -*-

// **********************************************************************
// *
// * legal mumbo jumbo
// *
// * (c) <year>, Cav
// * (utg v<utgversion>)
// ***********************************************************************
// File:   <filename>
// Author: <author>
/* About:  <description>
 *************************************************************************/

