<@header>
<@ifndef>

   `include "basic.sv"
// (`includes go here)

// class: <template>_c
// (Describe me)
class <template>_c extends base_test_c;
   `uvm_component_utils_begin(<template>_c)
   `uvm_component_utils_end

<@section_border>
   // Group: Configuration Fields

<@section_border>
   // Group: Fields

<@phases>
endclass : <template>_c

<@endif>
