<@header>
<@ifndef>

// `includes go here

// class: <class_name>
// (Describe me)
class <class_name> extends uvm_sequencer;
   `uvm_component_utils_begin(<vkit_name>_pkg::<class_name>)
   `uvm_component_utils_end

<@section_border>
   // Group: Configuration Fields

<@section_border>
   // Group: TLM Ports

<@section_border>
   // Group: Sequencer references
   // (put references to other sequencers here)

<@section_border>
   // Group: Fields

<@phases>
endclass : <class_name>


<@endif>
