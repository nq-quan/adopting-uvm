   ////////////////////////////////////////////
