<@header>
<@ifndef>
   
// (`includes go here)

// class: <name>_c
// (Describe me)
class <name>_c extends uvm_<template>;
   `uvm_component_utils_begin(<pkg_name>_pkg::<name>_c)
   `uvm_component_utils_end

<@section_border>
   // Group: Configuration Fields

<@section_border>
   // Group: TLM Ports
   
<@section_border>
   // Group: Fields

<@phases>
endclass : <name>_c
   
<@endif>
   