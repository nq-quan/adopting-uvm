<@header>

// (`includes of macros may go here)
`include "uvm_macros.svh"

// package: <class_name>
// (Describe me)
package <class_name>;

<@section_border>
   // Group: Imports
   import uvm_pkg::*;

<@section_border>
   // Group: Includes
   // (`include package member files here, alphabetically.)

endpackage : <class_name>


