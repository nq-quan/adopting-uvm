<@header>
<@ifndef>

// class: <class_name>
// (Describe me)
interface <class_name>(input logic clk, input logic rst_n);
   import uvm_pkg::*;

<@section_border>
   // Group: Signals

<@section_border>
   // Group: Clocking blocks

<@section_border>
   // Group: Modports

<@section_border>
   // Group: Methods

<@section_border>
   // Group: Assertions

endinterface : <class_name>

<@endif>
