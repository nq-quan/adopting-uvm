<@header>
<@ifndef>

// (`includes go here)

// class: <name>
// (Describe me)
class <class_name> extends uvm_<template>;
   `uvm_component_utils_begin(<vkit_name>_pkg::<name>)
   `uvm_component_utils_end

<@section_border>
   // Group: Configuration Fields

<@section_border>
   // Group: TLM Ports

<@section_border>
   // Group: Fields

<@phases>
endclass : <name>

<@endif>
