<@header>
<@ifndef>

   `include "base_test.sv"
// (`includes go here)

// class: <class_name>
// (Describe me)
class <class_name> extends base_test_c;
   `uvm_component_utils_begin(<class_name>)
   `uvm_component_utils_end

<@section_border>
   // Group: Configuration Fields

<@section_border>
   // Group: Fields

<@phases>
endclass : <class_name>

<@endif>
