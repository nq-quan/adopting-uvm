
// **********************************************************************
// *
// * legal mumbo jumbo
// *
// * (c) <year>
// * (utg v<utgversion>)
// ***********************************************************************
// File:   <filename>
// Author: <author>
/* About:  <description>
 *************************************************************************/

