<@header>
<@ifndef>

// `includes go here


<@endif>
         