//-*- mode: Verilog; verilog-indent-level: 3; indent-tabs-mode: nil; tab-width: 1 -*-

// **********************************************************************
// *
// * legal mumbo jumbo
// *
// * (c) 2012, Caviu
// * (utg v0.3.3)
// ***********************************************************************
// File:   cn_clk_mon.sv
// Author: jschroeder
/* About:  Clock Monitor

 *************************************************************************/

`ifndef __CN_CLK_MON_SV__
 `define __CN_CLK_MON_SV__

// Class: clock_mon_c
// A monitor for clocks that are generated by the DUT. Checks for correct
// period of the clock, whether the clock should be enabled or not, and checks
// that transitions are glitch-free.
//
// *extends <uvm_monitor>*
class clk_mon_c extends uvm_monitor;

   `uvm_component_utils_begin(cn_pkg::clk_mon_c)
      `uvm_field_string(intf_name,     UVM_ALL_ON)
      `uvm_field_int(max_period_ps,    UVM_ALL_ON)
      `uvm_field_int(initial_period_ps, UVM_ALL_ON)
      `uvm_field_int(disabled_state,   UVM_ALL_ON)
      `uvm_field_int(jitter_tolerance_pct, UVM_ALL_ON)
      `uvm_field_int(transition_timeout_ps, UVM_ALL_ON)
      `uvm_field_int(enable_checking,  UVM_ALL_ON)
      `uvm_field_int(auto_enable_checking, UVM_ALL_ON)
   `uvm_component_utils_end

   typedef struct {
      bit         valid;
      int         new_period_ps;
      realtime    transition_by;
   } transition_s;
   
   //--------------------------------------------------------------------------
   // Group: Configuration Fields

   // Field: intf_name
   // Name in the resource database under which the vintf is stored. The scope
   // under which it is stored is "cn_pkg::clk_intf".
   string intf_name = "clk_intf";

   // Field: max_period_ps
   // An upper bound on the period of the clock. If no transitions are seen in
   // this time interval, the clock is considered disabled.
   int    max_period_ps;

   // Field: initial_period_ps
   // The initial period of the clock when checking is started. A value of 0
   // means that the clock is expected to be disabled.
   int    initial_period_ps = 0;

   // Field: disabled_state
   // The expected state of the clock when it is disabled.
   bit    disabled_state = 0;
   
   // Field: jitter_tolerance_pct
   // Percentage variation allowed in the period of the clock while still
   // considering the period correct.
   int    jitter_tolerance_pct = 2;

   // Field: transition_timeout_ps
   // When the user indicates that the clock period will change, or that the
   // clock will be enabled or disabled, the change must happen within this
   // time period.
   int    transition_timeout_ps;

   // Field: enable_checking
   // Checking loop runs while enable_checking is 1.
   bit    enable_checking = 0;

   // Field: auto_enable_checking
   // Set to 0 to prevent checking from starting automatically in
   // pre_configure_phase.
   bit    auto_enable_checking = 1;
   
   //--------------------------------------------------------------------------
   // Group: Fields

   // interface to clock
   virtual cn_clk_intf clk_vi;

   // Last time we saw a clock edge. Used for calculating the half period.
   // Set to 0 when the clock is disabled.
   realtime last_clk_time = 0;
   
   // Bounds for the half period of the clock.
   realtime min_half_period;
   realtime max_half_period;

   // Flags that tell us if we've thrown certain errors. These are used to
   // avoid repeating ourselves.
   bit      clock_unknown_error = 0;
   bit      clock_transition_timeout_error = 0;
   bit      clock_period_error = 0;
   
   // Set by a call to <expect_transition>.
   transition_s next_transition;
   
   //--------------------------------------------------------------------------
   // Group: Methods

   ////////////////////////////////////////////
   // Constructor: new
   // Standard uvm_component constructor.
   function new(string name="clk_mon", uvm_component parent=null);
      super.new(name, parent);
   endfunction : new

   ////////////////////////////////////////////
   // Function: expect_transition
   // Expect a transition of the clock to a new period or for the clock
   // to be enabled or disabled.
   //
   // Arguments:
   //   new_period_ps - The new period of the clock in ps. A value of 0 means
   //     to expect the clock to be disabled.
   function void expect_transition(int new_period_ps);
      if (new_period_ps == 0 && last_clk_time == 0.0) begin
         `cn_warn(("Clock is already disabled"))
         return;
      end
      
      next_transition.valid = 1;
      next_transition.new_period_ps = new_period_ps;
      next_transition.transition_by = $realtime + transition_timeout_ps * 1ps;
   endfunction : expect_transition
   
   ////////////////////////////////////////////
   // Function: build_phase
   // Hook up to the virtual interface.
   virtual function void build_phase(uvm_phase phase);
      super.build_phase(phase);

      // get the interface
      `cn_get_intf(virtual cn_clk_intf, "cn_pkg::clk_intf", intf_name, clk_vi)

   endfunction : build_phase
   
   ////////////////////////////////////////////
   // Start checking in pre_configure_phase.
   virtual task pre_configure_phase(uvm_phase phase);
      super.pre_configure_phase(phase);
      if (auto_enable_checking) begin
         enable_checking = 1;
      end
   endtask : pre_configure_phase
   
   ////////////////////////////////////////////
   // Function: run_phase
   // Monitor the clock.
   virtual task run_phase(uvm_phase phase);

      forever begin
         wait (enable_checking == 1);

         // Force to disabled state.
         last_clk_time = 0.0;
         clock_transition_timeout_error = 0;
         clock_period_error = 0;

         // If starting in the disabled state, make sure the clock is in the
         // proper state.
         if (initial_period_ps == 0) begin
            if (clk_vi.clk !== disabled_state) begin
               `cn_err(("Clock is disabled, but is in the wrong state at initialization."))
            end
         end

         // If starting in the enabled state, set things to look like we're
         // transitioning from a disabled state. This works cleanly with the
         // main checking loop.
         else begin
            expect_transition(initial_period_ps);
         end

         while (enable_checking) begin
            logic last_clk;
         
            // Wait for either the next clock edge, or a maximum timeout period.
            last_clk = clk_vi.clk;
            fork
               wait (! enable_checking);
               #(max_period_ps * 1ps);
               @(clk_vi.clk);
            join_any
            disable fork;

            if (! enable_checking) begin
               continue;
            end
            
            // If clock is unknown, this is an error.
            if ($isunknown(clk_vi.clk)) begin
               if (! clock_unknown_error) begin
                  `cn_err(("Clock is unknown"))
               end
               clock_unknown_error = 1;
            end
            else begin
               clock_unknown_error = 0;
            end

            // If we saw an edge, the clock is running.
            if (clk_vi.clk !== last_clk) begin

               // If transitioning from a disabled state, make sure we're
               // expecting a transition.
               if (last_clk_time == 0.0) begin
                  if (! next_transition.valid) begin
                     `cn_err(("Saw a clock edge while clock should be disabled."))
                  end

                  // Calculate the new expected period.
                  else begin
                     `cn_dbg(UVM_MEDIUM, ("Clock %0s went from inactive to active with period %0d ps",
                                          intf_name,
                                          next_transition.new_period_ps))
                  
                     min_half_period = next_transition.new_period_ps * 1ps / 2.0 * (100.0 - jitter_tolerance_pct) / 100.0;
                     max_half_period = next_transition.new_period_ps * 1ps / 2.0 * (100.0 + jitter_tolerance_pct) / 100.0;
                     next_transition.valid = 0;
                     clock_period_error = 0;
                     clock_transition_timeout_error = 0;
                  end
               end

               // If not transitioning from a disbled state, calculate the half
               // period that was observed.
               else begin
                  realtime half_period_width;
            
                  half_period_width = $realtime - last_clk_time;

                  // If we're expecting a transition to a different period (not
                  // to a disabled clock), check if we've transitioned.
                  if (next_transition.valid && next_transition.new_period_ps != 0) begin

                     // Make sure we don't time out waiting for the transition.
                     if ($realtime > next_transition.transition_by) begin
                        if (! clock_transition_timeout_error) begin
                           `cn_err(("Clock did not transition to new period in the allotted time."))
                        end
                        clock_transition_timeout_error = 1;
                     end

                     // Check for clock glitches during the transition. A glitch
                     // is a half period that is less than both the old or new
                     // half periods.
                     if (half_period_width < min_half_period &&
                         half_period_width < next_transition.new_period_ps * 1ps / 2 * (100 - jitter_tolerance_pct) / 100) begin

                        `cn_err(("Clock glitched"))
                     end

                     // Check if the clock switched to the new period. It is
                     // considered switched if either the half period does not
                     // fit the old half period or it does fit the new half
                     // period. (The second clause covers the improbable case of
                     // old and new half period ranges that overlap.)
                     if (! (half_period_width inside {[min_half_period:max_half_period]} ||
                            half_period_width inside {[next_transition.new_period_ps * 1ps / 2 * (100 - jitter_tolerance_pct) / 100:
                                                       next_transition.new_period_ps * 1ps / 2 * (100 + jitter_tolerance_pct) / 100]})) begin
                     
                        `cn_dbg(UVM_MEDIUM, ("Clock %0s changed period to %0d ps",
                                             intf_name,
                                             next_transition.new_period_ps))
                     
                        min_half_period = next_transition.new_period_ps * 1ps / 2 * (100 - jitter_tolerance_pct) / 100;
                        max_half_period = next_transition.new_period_ps * 1ps / 2 * (100 + jitter_tolerance_pct) / 100;
                        next_transition.valid = 0;
                        clock_period_error = 0;
                        clock_transition_timeout_error = 0;
                     end
                  end

                  // If not expecting a transition, make sure the clock is the
                  // expected period.
                  else begin

                     // If we're expecting a transition to a disabled clock,
                     // check for timeout.
                     if (next_transition.valid && $realtime > next_transition.transition_by) begin
                        if (! clock_transition_timeout_error) begin
                           `cn_err(("Clock did not transition to new period in the allotted time."))
                        end
                        clock_transition_timeout_error = 1;
                     end

                     // Check the clock period.
                     if (! (half_period_width inside {[min_half_period:max_half_period]})) begin
                        if (! clock_period_error) begin
                           `cn_err(("Clock period is not as expected"))
                        end
                        clock_period_error = 1;
                     end
                  end
               end
            
               last_clk_time = $realtime;
            end

            // If we didn't see an edge, assume the clock is disabled.
            else begin

               // If transitioning from an enabled state, make sure we're
               // expecting a transition to a disabled state.
               if (last_clk_time != 0.0) begin
                  `cn_dbg(UVM_MEDIUM, ("Clock %0s went from active to inactive", intf_name))
               
                  if (! next_transition.valid || next_transition.new_period_ps != 0) begin
                     `cn_err(("Clock went inactive unexpectedly."))
                  end

                  if (clk_vi.clk !== disabled_state) begin
                     `cn_err(("Clock is disabled, but is in the wrong state"))
                  end
               
                  last_clk_time = 0;
                  next_transition.valid = 0;
                  clock_period_error = 0;
                  clock_transition_timeout_error = 0;
               end

               // If expecting a transition, check for timeout.
               if (next_transition.valid && $realtime > next_transition.transition_by) begin
                  if (! clock_transition_timeout_error) begin
                     `cn_err(("Clock did not transition to enabled state in the allotted time."))
                  end
                  clock_transition_timeout_error = 1;
               end
            end
         end
      end
   endtask : run_phase
   
endclass : clk_mon_c

`endif // __CN_CLK_MON_SV__