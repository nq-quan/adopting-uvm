<@header>
<@ifndef>

// class: <template>
// (Describe me)
interface <template>(input logic clk, input logic rst_n);

<@section_border>
   // Group: Signals

<@section_border>
   // Group: Clocking blocks

<@section_border>
   // Group: Modports

<@section_border>
   // Group: Methods

<@section_border>
   // Group: Assertions

endinterface : <template>

<@endif>
