//****************************************************************************************
