<@header>
<@ifndef>
   
// (`includes go here)

// (your first sequence!)
<@vseq>

<@endif>
   