`ifndef __<FILENAME>_SV__
   `define __<FILENAME>_SV__

<?selftest>
    `include "cn_self_test.sv"
<?end>
