
// **********************************************************************
// *
// * legal mumbo jumbo
// *
// * (c) 2013
// * (utg v0.10)
// ***********************************************************************
// File:   res_types.sv
// Author: bhunter
/* About:  Types file.
 *************************************************************************/

`ifndef __RES_TYPES_SV__
   `define __RES_TYPES_SV__

typedef bit[31:0]  result_t;


`endif // __RES_TYPES_SV__
