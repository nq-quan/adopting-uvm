<@header>

// (`includes of macros may go here)
`include "uvm_macros.svh"

// package: <pkg_name>_<template>
// (Describe me)
package <pkg_name>_<template>;

<@section_border>
   // Group: Imports
   import uvm_pkg::*;

<@section_border>
   // Group: Includes
   // (`include package member files here, alphabetically.)
   
endpackage : <pkg_name>_<template>
   

