   //----------------------------------------------------------------------------------------
