<@header>
<@ifndef>
   
// `includes go here

// class: <template>_c
// (Describe me)
class <template>_c extends uvm_sequencer;
   `uvm_component_utils_begin(<pkg_name>_pkg::<template>_c)
   `uvm_component_utils_end

<@section_border>
   // Group: Configuration Fields

<@section_border>
   // Group: TLM Ports

<@section_border>
   // Group: Sequencer references
   // (put references to other sequencers here)

<@section_border>
   // Group: Fields

<@phases>
endclass : <template>_c
   

<@endif>
   