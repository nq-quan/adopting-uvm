
// **********************************************************************
// *
// * legal mumbo jumbo
// *
// * (c) <year>, Cav
// * (utg v<utgversion>)
// ***********************************************************************
// File:   <filename>
// Author: <author>
/* About:  <description>
 *************************************************************************/

