`ifndef __<FILENAME>_SV__
   `define __<FILENAME>_SV__
