<@header>
<@ifndef>

// (`includes go here)

// class: <class_name>
// (Describe me)
class drv_c extends uvm_driver#(<reqType>,<rspType>);
   `uvm_component_utils_begin(<vkit_name>_pkg::<class_name>)
   `uvm_component_utils_end

<@section_border>
   // Group: Configuration Fields

<@section_border>
   // Group: TLM Ports

<@section_border>
   // Group: Fields

<@phases>
endclass : <class_name>

<@endif>