`endif // __<FILENAME>_SV__
